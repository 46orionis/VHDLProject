  
VDS